module menu
